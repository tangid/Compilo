`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:44:02 05/03/2018 
// Design Name: 
// Module Name:    ual 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ual(
    input [15:0] A,
    input [15:0] B,
    input [4:0] op,
    output [15:0] S,
    output [4:0] flag
    );


endmodule
